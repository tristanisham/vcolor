module color

const (
	//Black sets text color to black
	Black = "30"
	//DarkRed sets text color to dark red
	DarkRed = "31"
	//DarkGreen sets text color to dark green
	DarkGreen = "32"
	//DarkYellow sets text color to dark yellow
	DarkYellow = "33"
	//DarkBlue sets text color to dark blue
	DarkBlue = "34"
	//DarkMagenta sets text color to dark magenta
	DarkMagenta = "35"
	//DarkCyan sets text color to dark cyan
	DarkCyan = "36"
	//LightGray sets text color to light gray
	LightGray = "37"
	//DarkGray sets text color to dark gray
	DarkGray = "90"
	//LightRed sets text color to light red
	LightRed = "91"
	//LightGreen sets text color to light green
	LightGreen = "92"
	//LightYellow sets text color to light yellow
	LightYellow = "93"
	//LightBlue sets text color to light blue
	LightBlue = "94"
	//LightMagenta sets text color to light magenta
	LightMagenta = "95"
	//LightCyan sets text color to light cyan
	LightCyan = "96"
	//White sets text color to White
	White = "97"

	BgBlack        = "40"
	BgDarkRed      = "41"
	BgDarkGreen    = "42"
	BgDarkYellow   = "43"
	BgDarkBlue     = "44"
	BgDarkCyan     = "46"
	BgLightGray    = "100"
	BgLightRed     = "101"
	BgLightGreen   = "102"
	BgLightYellow  = "103"
	BgLightBlue    = "104"
	BgLightMagenta = "105"
	BgLightCyan    = "106"
	BgWhite        = "107"
	//
	Bold        = "1"
	Underline   = "4"
	NoUnderline = "24"
	// ReverseText  = "7"
	PositiveText = "27"
	Reset        = "\033[0m"
)